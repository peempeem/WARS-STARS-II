// soc.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module soc (
		input  wire        clk_clk,          //        clk.clk
		input  wire        reset_reset_n,    //      reset.reset_n
		output wire        sdram_clk_clk,    //  sdram_clk.clk
		output wire [12:0] sdram_wire_addr,  // sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,    //           .ba
		output wire        sdram_wire_cas_n, //           .cas_n
		output wire        sdram_wire_cke,   //           .cke
		output wire        sdram_wire_cs_n,  //           .cs_n
		inout  wire [15:0] sdram_wire_dq,    //           .dq
		output wire [1:0]  sdram_wire_dqm,   //           .dqm
		output wire        sdram_wire_ras_n, //           .ras_n
		output wire        sdram_wire_we_n,  //           .we_n
		input  wire        spi0_MISO,        //       spi0.MISO
		output wire        spi0_MOSI,        //           .MOSI
		output wire        spi0_SCLK,        //           .SCLK
		output wire        spi0_SS_n,        //           .SS_n
		input  wire        usb_gpx_export,   //    usb_gpx.export
		input  wire        usb_irq_export,   //    usb_irq.export
		output wire        usb_rst_export,   //    usb_rst.export
		output wire [3:0]  vga_port_blue,    //   vga_port.blue
		output wire [3:0]  vga_port_green,   //           .green
		output wire        vga_port_hs,      //           .hs
		output wire [3:0]  vga_port_red,     //           .red
		output wire        vga_port_vs       //           .vs
	);

	wire         pll_c0_clk;                                                       // pll:c0 -> [mm_interconnect_0:pll_c0_clk, rst_controller_002:clk, sdram:clk]
	wire         pll_c2_clk;                                                       // pll:c2 -> [graphics_drawing_unit_0:clk1, mm_interconnect_0:pll_c2_clk, rst_controller_003:clk]
	wire         pll_c3_clk;                                                       // pll:c3 -> Timer_64Bit_0:clk1
	wire  [31:0] vga_display_0_avalon_master_readdata;                             // mm_interconnect_0:vga_display_0_avalon_master_readdata -> vga_display_0:avalon_master_readdata
	wire         vga_display_0_avalon_master_waitrequest;                          // mm_interconnect_0:vga_display_0_avalon_master_waitrequest -> vga_display_0:avalon_master_waitrequest
	wire         vga_display_0_avalon_master_read;                                 // vga_display_0:avalon_master_read -> mm_interconnect_0:vga_display_0_avalon_master_read
	wire  [31:0] vga_display_0_avalon_master_address;                              // vga_display_0:avalon_master_address -> mm_interconnect_0:vga_display_0_avalon_master_address
	wire         vga_display_0_avalon_master_readdatavalid;                        // mm_interconnect_0:vga_display_0_avalon_master_readdatavalid -> vga_display_0:avalon_master_readdatavalid
	wire   [4:0] vga_display_0_avalon_master_burstcount;                           // vga_display_0:avalon_master_burstcount -> mm_interconnect_0:vga_display_0_avalon_master_burstcount
	wire  [31:0] graphics_drawing_unit_0_avalon_master_readdata;                   // mm_interconnect_0:graphics_drawing_unit_0_avalon_master_readdata -> graphics_drawing_unit_0:avalon_master_readdata
	wire         graphics_drawing_unit_0_avalon_master_waitrequest;                // mm_interconnect_0:graphics_drawing_unit_0_avalon_master_waitrequest -> graphics_drawing_unit_0:avalon_master_waitrequest
	wire  [31:0] graphics_drawing_unit_0_avalon_master_address;                    // graphics_drawing_unit_0:avalon_master_address -> mm_interconnect_0:graphics_drawing_unit_0_avalon_master_address
	wire         graphics_drawing_unit_0_avalon_master_read;                       // graphics_drawing_unit_0:avalon_master_read -> mm_interconnect_0:graphics_drawing_unit_0_avalon_master_read
	wire   [3:0] graphics_drawing_unit_0_avalon_master_byteenable;                 // graphics_drawing_unit_0:avalon_master_byteenable -> mm_interconnect_0:graphics_drawing_unit_0_avalon_master_byteenable
	wire         graphics_drawing_unit_0_avalon_master_readdatavalid;              // mm_interconnect_0:graphics_drawing_unit_0_avalon_master_readdatavalid -> graphics_drawing_unit_0:avalon_master_readdatavalid
	wire   [1:0] graphics_drawing_unit_0_avalon_master_response;                   // mm_interconnect_0:graphics_drawing_unit_0_avalon_master_response -> graphics_drawing_unit_0:avalon_master_response
	wire  [31:0] graphics_drawing_unit_0_avalon_master_writedata;                  // graphics_drawing_unit_0:avalon_master_writedata -> mm_interconnect_0:graphics_drawing_unit_0_avalon_master_writedata
	wire         graphics_drawing_unit_0_avalon_master_write;                      // graphics_drawing_unit_0:avalon_master_write -> mm_interconnect_0:graphics_drawing_unit_0_avalon_master_write
	wire         graphics_drawing_unit_0_avalon_master_writeresponsevalid;         // mm_interconnect_0:graphics_drawing_unit_0_avalon_master_writeresponsevalid -> graphics_drawing_unit_0:avalon_master_writeresponsevalid
	wire   [3:0] graphics_drawing_unit_0_avalon_master_burstcount;                 // graphics_drawing_unit_0:avalon_master_burstcount -> mm_interconnect_0:graphics_drawing_unit_0_avalon_master_burstcount
	wire  [31:0] nios2_gen2_0_data_master_readdata;                                // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                             // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                             // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [27:0] nios2_gen2_0_data_master_address;                                 // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                              // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                    // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                                   // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                               // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                         // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                      // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [27:0] nios2_gen2_0_instruction_master_address;                          // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                             // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_sdram_s1_chipselect;                            // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                              // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                           // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                               // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                  // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                            // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                         // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                 // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                             // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;         // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;      // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;          // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;             // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;            // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_vga_display_0_avalon_slave_readdata;            // vga_display_0:avalon_slave_readdata -> mm_interconnect_0:vga_display_0_avalon_slave_readdata
	wire   [2:0] mm_interconnect_0_vga_display_0_avalon_slave_address;             // mm_interconnect_0:vga_display_0_avalon_slave_address -> vga_display_0:avalon_slave_address
	wire         mm_interconnect_0_vga_display_0_avalon_slave_read;                // mm_interconnect_0:vga_display_0_avalon_slave_read -> vga_display_0:avalon_slave_read
	wire         mm_interconnect_0_vga_display_0_avalon_slave_write;               // mm_interconnect_0:vga_display_0_avalon_slave_write -> vga_display_0:avalon_slave_write
	wire  [31:0] mm_interconnect_0_vga_display_0_avalon_slave_writedata;           // mm_interconnect_0:vga_display_0_avalon_slave_writedata -> vga_display_0:avalon_slave_writedata
	wire  [31:0] mm_interconnect_0_graphics_drawing_unit_0_avalon_slave_readdata;  // graphics_drawing_unit_0:avalon_slave_readdata -> mm_interconnect_0:graphics_drawing_unit_0_avalon_slave_readdata
	wire  [10:0] mm_interconnect_0_graphics_drawing_unit_0_avalon_slave_address;   // mm_interconnect_0:graphics_drawing_unit_0_avalon_slave_address -> graphics_drawing_unit_0:avalon_slave_address
	wire         mm_interconnect_0_graphics_drawing_unit_0_avalon_slave_read;      // mm_interconnect_0:graphics_drawing_unit_0_avalon_slave_read -> graphics_drawing_unit_0:avalon_slave_read
	wire         mm_interconnect_0_graphics_drawing_unit_0_avalon_slave_write;     // mm_interconnect_0:graphics_drawing_unit_0_avalon_slave_write -> graphics_drawing_unit_0:avalon_slave_write
	wire  [31:0] mm_interconnect_0_graphics_drawing_unit_0_avalon_slave_writedata; // mm_interconnect_0:graphics_drawing_unit_0_avalon_slave_writedata -> graphics_drawing_unit_0:avalon_slave_writedata
	wire  [31:0] mm_interconnect_0_timer_64bit_0_avalon_slave_readdata;            // Timer_64Bit_0:avalon_slave_readdata -> mm_interconnect_0:Timer_64Bit_0_avalon_slave_readdata
	wire   [1:0] mm_interconnect_0_timer_64bit_0_avalon_slave_address;             // mm_interconnect_0:Timer_64Bit_0_avalon_slave_address -> Timer_64Bit_0:avalon_slave_address
	wire         mm_interconnect_0_timer_64bit_0_avalon_slave_read;                // mm_interconnect_0:Timer_64Bit_0_avalon_slave_read -> Timer_64Bit_0:avalon_slave_read
	wire         mm_interconnect_0_timer_64bit_0_avalon_slave_write;               // mm_interconnect_0:Timer_64Bit_0_avalon_slave_write -> Timer_64Bit_0:avalon_slave_write
	wire  [31:0] mm_interconnect_0_timer_64bit_0_avalon_slave_writedata;           // mm_interconnect_0:Timer_64Bit_0_avalon_slave_writedata -> Timer_64Bit_0:avalon_slave_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;            // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;             // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;          // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;       // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;           // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;              // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;             // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_pll_pll_slave_readdata;                         // pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_pll_pll_slave_address;                          // mm_interconnect_0:pll_pll_slave_address -> pll:address
	wire         mm_interconnect_0_pll_pll_slave_read;                             // mm_interconnect_0:pll_pll_slave_read -> pll:read
	wire         mm_interconnect_0_pll_pll_slave_write;                            // mm_interconnect_0:pll_pll_slave_write -> pll:write
	wire  [31:0] mm_interconnect_0_pll_pll_slave_writedata;                        // mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	wire  [31:0] mm_interconnect_0_usb_irq_s1_readdata;                            // usb_irq:readdata -> mm_interconnect_0:usb_irq_s1_readdata
	wire   [1:0] mm_interconnect_0_usb_irq_s1_address;                             // mm_interconnect_0:usb_irq_s1_address -> usb_irq:address
	wire  [31:0] mm_interconnect_0_usb_gpx_s1_readdata;                            // usb_gpx:readdata -> mm_interconnect_0:usb_gpx_s1_readdata
	wire   [1:0] mm_interconnect_0_usb_gpx_s1_address;                             // mm_interconnect_0:usb_gpx_s1_address -> usb_gpx:address
	wire         mm_interconnect_0_usb_rst_s1_chipselect;                          // mm_interconnect_0:usb_rst_s1_chipselect -> usb_rst:chipselect
	wire  [31:0] mm_interconnect_0_usb_rst_s1_readdata;                            // usb_rst:readdata -> mm_interconnect_0:usb_rst_s1_readdata
	wire   [1:0] mm_interconnect_0_usb_rst_s1_address;                             // mm_interconnect_0:usb_rst_s1_address -> usb_rst:address
	wire         mm_interconnect_0_usb_rst_s1_write;                               // mm_interconnect_0:usb_rst_s1_write -> usb_rst:write_n
	wire  [31:0] mm_interconnect_0_usb_rst_s1_writedata;                           // mm_interconnect_0:usb_rst_s1_writedata -> usb_rst:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                          // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                            // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [3:0] mm_interconnect_0_timer_0_s1_address;                             // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                               // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                           // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                 // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                   // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [9:0] mm_interconnect_0_onchip_memory2_0_s1_address;                    // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                 // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                      // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                  // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                      // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_spi_0_spi_control_port_chipselect;              // mm_interconnect_0:spi_0_spi_control_port_chipselect -> spi_0:spi_select
	wire  [15:0] mm_interconnect_0_spi_0_spi_control_port_readdata;                // spi_0:data_to_cpu -> mm_interconnect_0:spi_0_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_0_spi_control_port_address;                 // mm_interconnect_0:spi_0_spi_control_port_address -> spi_0:mem_addr
	wire         mm_interconnect_0_spi_0_spi_control_port_read;                    // mm_interconnect_0:spi_0_spi_control_port_read -> spi_0:read_n
	wire         mm_interconnect_0_spi_0_spi_control_port_write;                   // mm_interconnect_0:spi_0_spi_control_port_write -> spi_0:write_n
	wire  [15:0] mm_interconnect_0_spi_0_spi_control_port_writedata;               // mm_interconnect_0:spi_0_spi_control_port_writedata -> spi_0:data_from_cpu
	wire         irq_mapper_receiver0_irq;                                         // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                         // timer_0:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                         // spi_0:irq -> irq_mapper:receiver2_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                             // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                                   // rst_controller:reset_out -> [Timer_64Bit_0:reset, graphics_drawing_unit_0:reset, irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                               // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                               // rst_controller_001:reset_out -> [jtag_uart_0:rst_n, mm_interconnect_0:vga_display_0_reset_reset_bridge_in_reset_reset, pll:reset, spi_0:reset_n, sysid_qsys_0:reset_n, timer_0:reset_n, usb_gpx:reset_n, usb_irq:reset_n, usb_rst:reset_n, vga_display_0:reset]
	wire         nios2_gen2_0_debug_reset_request_reset;                           // nios2_gen2_0:debug_reset_request -> [rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_002_reset_out_reset;                               // rst_controller_002:reset_out -> [mm_interconnect_0:sdram_reset_reset_bridge_in_reset_reset, sdram:reset_n]
	wire         rst_controller_003_reset_out_reset;                               // rst_controller_003:reset_out -> mm_interconnect_0:graphics_drawing_unit_0_reset_reset_bridge_in_reset_reset

	Timer timer_64bit_0 (
		.reset                  (rst_controller_reset_out_reset),                         //        reset.reset
		.avalon_slave_address   (mm_interconnect_0_timer_64bit_0_avalon_slave_address),   // avalon_slave.address
		.avalon_slave_read      (mm_interconnect_0_timer_64bit_0_avalon_slave_read),      //             .read
		.avalon_slave_readdata  (mm_interconnect_0_timer_64bit_0_avalon_slave_readdata),  //             .readdata
		.avalon_slave_write     (mm_interconnect_0_timer_64bit_0_avalon_slave_write),     //             .write
		.avalon_slave_writedata (mm_interconnect_0_timer_64bit_0_avalon_slave_writedata), //             .writedata
		.clk1                   (pll_c3_clk),                                             //         clk1.clk
		.clk0                   (clk_clk)                                                 //         clk0.clk
	);

	graphics_drawing_unit graphics_drawing_unit_0 (
		.reset                            (rst_controller_reset_out_reset),                                   //         reset.reset
		.avalon_master_address            (graphics_drawing_unit_0_avalon_master_address),                    // avalon_master.address
		.avalon_master_burstcount         (graphics_drawing_unit_0_avalon_master_burstcount),                 //              .burstcount
		.avalon_master_read               (graphics_drawing_unit_0_avalon_master_read),                       //              .read
		.avalon_master_readdata           (graphics_drawing_unit_0_avalon_master_readdata),                   //              .readdata
		.avalon_master_waitrequest        (graphics_drawing_unit_0_avalon_master_waitrequest),                //              .waitrequest
		.avalon_master_writedata          (graphics_drawing_unit_0_avalon_master_writedata),                  //              .writedata
		.avalon_master_write              (graphics_drawing_unit_0_avalon_master_write),                      //              .write
		.avalon_master_byteenable         (graphics_drawing_unit_0_avalon_master_byteenable),                 //              .byteenable
		.avalon_master_readdatavalid      (graphics_drawing_unit_0_avalon_master_readdatavalid),              //              .readdatavalid
		.avalon_master_writeresponsevalid (graphics_drawing_unit_0_avalon_master_writeresponsevalid),         //              .writeresponsevalid
		.avalon_master_response           (graphics_drawing_unit_0_avalon_master_response),                   //              .response
		.avalon_slave_address             (mm_interconnect_0_graphics_drawing_unit_0_avalon_slave_address),   //  avalon_slave.address
		.avalon_slave_read                (mm_interconnect_0_graphics_drawing_unit_0_avalon_slave_read),      //              .read
		.avalon_slave_readdata            (mm_interconnect_0_graphics_drawing_unit_0_avalon_slave_readdata),  //              .readdata
		.avalon_slave_write               (mm_interconnect_0_graphics_drawing_unit_0_avalon_slave_write),     //              .write
		.avalon_slave_writedata           (mm_interconnect_0_graphics_drawing_unit_0_avalon_slave_writedata), //              .writedata
		.clk1                             (pll_c2_clk),                                                       //          clk1.clk
		.clk0                             (clk_clk)                                                           //          clk0.clk
	);

	soc_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	soc_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	soc_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	soc_pll pll (
		.clk                (clk_clk),                                   //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),        // inclk_interface_reset.reset
		.read               (mm_interconnect_0_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_pll_pll_slave_writedata), //                      .writedata
		.c0                 (pll_c0_clk),                                //                    c0.clk
		.c1                 (sdram_clk_clk),                             //                    c1.clk
		.c2                 (pll_c2_clk),                                //                    c2.clk
		.c3                 (pll_c3_clk),                                //                    c3.clk
		.scandone           (),                                          //           (terminated)
		.scandataout        (),                                          //           (terminated)
		.c4                 (),                                          //           (terminated)
		.areset             (1'b0),                                      //           (terminated)
		.locked             (),                                          //           (terminated)
		.phasedone          (),                                          //           (terminated)
		.phasecounterselect (3'b000),                                    //           (terminated)
		.phaseupdown        (1'b0),                                      //           (terminated)
		.phasestep          (1'b0),                                      //           (terminated)
		.scanclk            (1'b0),                                      //           (terminated)
		.scanclkena         (1'b0),                                      //           (terminated)
		.scandata           (1'b0),                                      //           (terminated)
		.configupdate       (1'b0)                                       //           (terminated)
	);

	soc_sdram sdram (
		.clk            (pll_c0_clk),                               //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	soc_spi_0 spi_0 (
		.clk           (clk_clk),                                             //              clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                 //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_0_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_0_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_0_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_0_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_0_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_0_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver2_irq),                            //              irq.irq
		.MISO          (spi0_MISO),                                           //         external.export
		.MOSI          (spi0_MOSI),                                           //                 .export
		.SCLK          (spi0_SCLK),                                           //                 .export
		.SS_n          (spi0_SS_n)                                            //                 .export
	);

	soc_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	soc_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	soc_usb_gpx usb_gpx (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_usb_gpx_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_usb_gpx_s1_readdata), //                    .readdata
		.in_port  (usb_gpx_export)                         // external_connection.export
	);

	soc_usb_gpx usb_irq (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_usb_irq_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_usb_irq_s1_readdata), //                    .readdata
		.in_port  (usb_irq_export)                         // external_connection.export
	);

	soc_usb_rst usb_rst (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_usb_rst_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_usb_rst_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_usb_rst_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_usb_rst_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_usb_rst_s1_readdata),   //                    .readdata
		.out_port   (usb_rst_export)                           // external_connection.export
	);

	vga_display vga_display_0 (
		.clk                         (clk_clk),                                                //         clock.clk
		.reset                       (rst_controller_001_reset_out_reset),                     //         reset.reset
		.blue                        (vga_port_blue),                                          //      vga_port.blue
		.green                       (vga_port_green),                                         //              .green
		.hs                          (vga_port_hs),                                            //              .hs
		.red                         (vga_port_red),                                           //              .red
		.vs                          (vga_port_vs),                                            //              .vs
		.avalon_master_read          (vga_display_0_avalon_master_read),                       // avalon_master.read
		.avalon_master_readdata      (vga_display_0_avalon_master_readdata),                   //              .readdata
		.avalon_master_readdatavalid (vga_display_0_avalon_master_readdatavalid),              //              .readdatavalid
		.avalon_master_waitrequest   (vga_display_0_avalon_master_waitrequest),                //              .waitrequest
		.avalon_master_address       (vga_display_0_avalon_master_address),                    //              .address
		.avalon_master_burstcount    (vga_display_0_avalon_master_burstcount),                 //              .burstcount
		.avalon_slave_address        (mm_interconnect_0_vga_display_0_avalon_slave_address),   //  avalon_slave.address
		.avalon_slave_read           (mm_interconnect_0_vga_display_0_avalon_slave_read),      //              .read
		.avalon_slave_write          (mm_interconnect_0_vga_display_0_avalon_slave_write),     //              .write
		.avalon_slave_readdata       (mm_interconnect_0_vga_display_0_avalon_slave_readdata),  //              .readdata
		.avalon_slave_writedata      (mm_interconnect_0_vga_display_0_avalon_slave_writedata)  //              .writedata
	);

	soc_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                             (clk_clk),                                                          //                                           clk_0_clk.clk
		.pll_c0_clk                                                (pll_c0_clk),                                                       //                                              pll_c0.clk
		.pll_c2_clk                                                (pll_c2_clk),                                                       //                                              pll_c2.clk
		.graphics_drawing_unit_0_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                               // graphics_drawing_unit_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset            (rst_controller_reset_out_reset),                                   //            nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.sdram_reset_reset_bridge_in_reset_reset                   (rst_controller_002_reset_out_reset),                               //                   sdram_reset_reset_bridge_in_reset.reset
		.vga_display_0_reset_reset_bridge_in_reset_reset           (rst_controller_001_reset_out_reset),                               //           vga_display_0_reset_reset_bridge_in_reset.reset
		.graphics_drawing_unit_0_avalon_master_address             (graphics_drawing_unit_0_avalon_master_address),                    //               graphics_drawing_unit_0_avalon_master.address
		.graphics_drawing_unit_0_avalon_master_waitrequest         (graphics_drawing_unit_0_avalon_master_waitrequest),                //                                                    .waitrequest
		.graphics_drawing_unit_0_avalon_master_burstcount          (graphics_drawing_unit_0_avalon_master_burstcount),                 //                                                    .burstcount
		.graphics_drawing_unit_0_avalon_master_byteenable          (graphics_drawing_unit_0_avalon_master_byteenable),                 //                                                    .byteenable
		.graphics_drawing_unit_0_avalon_master_read                (graphics_drawing_unit_0_avalon_master_read),                       //                                                    .read
		.graphics_drawing_unit_0_avalon_master_readdata            (graphics_drawing_unit_0_avalon_master_readdata),                   //                                                    .readdata
		.graphics_drawing_unit_0_avalon_master_readdatavalid       (graphics_drawing_unit_0_avalon_master_readdatavalid),              //                                                    .readdatavalid
		.graphics_drawing_unit_0_avalon_master_write               (graphics_drawing_unit_0_avalon_master_write),                      //                                                    .write
		.graphics_drawing_unit_0_avalon_master_writedata           (graphics_drawing_unit_0_avalon_master_writedata),                  //                                                    .writedata
		.graphics_drawing_unit_0_avalon_master_response            (graphics_drawing_unit_0_avalon_master_response),                   //                                                    .response
		.graphics_drawing_unit_0_avalon_master_writeresponsevalid  (graphics_drawing_unit_0_avalon_master_writeresponsevalid),         //                                                    .writeresponsevalid
		.nios2_gen2_0_data_master_address                          (nios2_gen2_0_data_master_address),                                 //                            nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                      (nios2_gen2_0_data_master_waitrequest),                             //                                                    .waitrequest
		.nios2_gen2_0_data_master_byteenable                       (nios2_gen2_0_data_master_byteenable),                              //                                                    .byteenable
		.nios2_gen2_0_data_master_read                             (nios2_gen2_0_data_master_read),                                    //                                                    .read
		.nios2_gen2_0_data_master_readdata                         (nios2_gen2_0_data_master_readdata),                                //                                                    .readdata
		.nios2_gen2_0_data_master_write                            (nios2_gen2_0_data_master_write),                                   //                                                    .write
		.nios2_gen2_0_data_master_writedata                        (nios2_gen2_0_data_master_writedata),                               //                                                    .writedata
		.nios2_gen2_0_data_master_debugaccess                      (nios2_gen2_0_data_master_debugaccess),                             //                                                    .debugaccess
		.nios2_gen2_0_instruction_master_address                   (nios2_gen2_0_instruction_master_address),                          //                     nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest               (nios2_gen2_0_instruction_master_waitrequest),                      //                                                    .waitrequest
		.nios2_gen2_0_instruction_master_read                      (nios2_gen2_0_instruction_master_read),                             //                                                    .read
		.nios2_gen2_0_instruction_master_readdata                  (nios2_gen2_0_instruction_master_readdata),                         //                                                    .readdata
		.vga_display_0_avalon_master_address                       (vga_display_0_avalon_master_address),                              //                         vga_display_0_avalon_master.address
		.vga_display_0_avalon_master_waitrequest                   (vga_display_0_avalon_master_waitrequest),                          //                                                    .waitrequest
		.vga_display_0_avalon_master_burstcount                    (vga_display_0_avalon_master_burstcount),                           //                                                    .burstcount
		.vga_display_0_avalon_master_read                          (vga_display_0_avalon_master_read),                                 //                                                    .read
		.vga_display_0_avalon_master_readdata                      (vga_display_0_avalon_master_readdata),                             //                                                    .readdata
		.vga_display_0_avalon_master_readdatavalid                 (vga_display_0_avalon_master_readdatavalid),                        //                                                    .readdatavalid
		.graphics_drawing_unit_0_avalon_slave_address              (mm_interconnect_0_graphics_drawing_unit_0_avalon_slave_address),   //                graphics_drawing_unit_0_avalon_slave.address
		.graphics_drawing_unit_0_avalon_slave_write                (mm_interconnect_0_graphics_drawing_unit_0_avalon_slave_write),     //                                                    .write
		.graphics_drawing_unit_0_avalon_slave_read                 (mm_interconnect_0_graphics_drawing_unit_0_avalon_slave_read),      //                                                    .read
		.graphics_drawing_unit_0_avalon_slave_readdata             (mm_interconnect_0_graphics_drawing_unit_0_avalon_slave_readdata),  //                                                    .readdata
		.graphics_drawing_unit_0_avalon_slave_writedata            (mm_interconnect_0_graphics_drawing_unit_0_avalon_slave_writedata), //                                                    .writedata
		.jtag_uart_0_avalon_jtag_slave_address                     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),          //                       jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),            //                                                    .write
		.jtag_uart_0_avalon_jtag_slave_read                        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),             //                                                    .read
		.jtag_uart_0_avalon_jtag_slave_readdata                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),         //                                                    .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),        //                                                    .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                 (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),      //                                                    .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),       //                                                    .chipselect
		.nios2_gen2_0_debug_mem_slave_address                      (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),           //                        nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),             //                                                    .write
		.nios2_gen2_0_debug_mem_slave_read                         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),              //                                                    .read
		.nios2_gen2_0_debug_mem_slave_readdata                     (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),          //                                                    .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                    (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),         //                                                    .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),        //                                                    .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                  (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),       //                                                    .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                  (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),       //                                                    .debugaccess
		.onchip_memory2_0_s1_address                               (mm_interconnect_0_onchip_memory2_0_s1_address),                    //                                 onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                 (mm_interconnect_0_onchip_memory2_0_s1_write),                      //                                                    .write
		.onchip_memory2_0_s1_readdata                              (mm_interconnect_0_onchip_memory2_0_s1_readdata),                   //                                                    .readdata
		.onchip_memory2_0_s1_writedata                             (mm_interconnect_0_onchip_memory2_0_s1_writedata),                  //                                                    .writedata
		.onchip_memory2_0_s1_byteenable                            (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                 //                                                    .byteenable
		.onchip_memory2_0_s1_chipselect                            (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                 //                                                    .chipselect
		.onchip_memory2_0_s1_clken                                 (mm_interconnect_0_onchip_memory2_0_s1_clken),                      //                                                    .clken
		.pll_pll_slave_address                                     (mm_interconnect_0_pll_pll_slave_address),                          //                                       pll_pll_slave.address
		.pll_pll_slave_write                                       (mm_interconnect_0_pll_pll_slave_write),                            //                                                    .write
		.pll_pll_slave_read                                        (mm_interconnect_0_pll_pll_slave_read),                             //                                                    .read
		.pll_pll_slave_readdata                                    (mm_interconnect_0_pll_pll_slave_readdata),                         //                                                    .readdata
		.pll_pll_slave_writedata                                   (mm_interconnect_0_pll_pll_slave_writedata),                        //                                                    .writedata
		.sdram_s1_address                                          (mm_interconnect_0_sdram_s1_address),                               //                                            sdram_s1.address
		.sdram_s1_write                                            (mm_interconnect_0_sdram_s1_write),                                 //                                                    .write
		.sdram_s1_read                                             (mm_interconnect_0_sdram_s1_read),                                  //                                                    .read
		.sdram_s1_readdata                                         (mm_interconnect_0_sdram_s1_readdata),                              //                                                    .readdata
		.sdram_s1_writedata                                        (mm_interconnect_0_sdram_s1_writedata),                             //                                                    .writedata
		.sdram_s1_byteenable                                       (mm_interconnect_0_sdram_s1_byteenable),                            //                                                    .byteenable
		.sdram_s1_readdatavalid                                    (mm_interconnect_0_sdram_s1_readdatavalid),                         //                                                    .readdatavalid
		.sdram_s1_waitrequest                                      (mm_interconnect_0_sdram_s1_waitrequest),                           //                                                    .waitrequest
		.sdram_s1_chipselect                                       (mm_interconnect_0_sdram_s1_chipselect),                            //                                                    .chipselect
		.spi_0_spi_control_port_address                            (mm_interconnect_0_spi_0_spi_control_port_address),                 //                              spi_0_spi_control_port.address
		.spi_0_spi_control_port_write                              (mm_interconnect_0_spi_0_spi_control_port_write),                   //                                                    .write
		.spi_0_spi_control_port_read                               (mm_interconnect_0_spi_0_spi_control_port_read),                    //                                                    .read
		.spi_0_spi_control_port_readdata                           (mm_interconnect_0_spi_0_spi_control_port_readdata),                //                                                    .readdata
		.spi_0_spi_control_port_writedata                          (mm_interconnect_0_spi_0_spi_control_port_writedata),               //                                                    .writedata
		.spi_0_spi_control_port_chipselect                         (mm_interconnect_0_spi_0_spi_control_port_chipselect),              //                                                    .chipselect
		.sysid_qsys_0_control_slave_address                        (mm_interconnect_0_sysid_qsys_0_control_slave_address),             //                          sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                       (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),            //                                                    .readdata
		.timer_0_s1_address                                        (mm_interconnect_0_timer_0_s1_address),                             //                                          timer_0_s1.address
		.timer_0_s1_write                                          (mm_interconnect_0_timer_0_s1_write),                               //                                                    .write
		.timer_0_s1_readdata                                       (mm_interconnect_0_timer_0_s1_readdata),                            //                                                    .readdata
		.timer_0_s1_writedata                                      (mm_interconnect_0_timer_0_s1_writedata),                           //                                                    .writedata
		.timer_0_s1_chipselect                                     (mm_interconnect_0_timer_0_s1_chipselect),                          //                                                    .chipselect
		.Timer_64Bit_0_avalon_slave_address                        (mm_interconnect_0_timer_64bit_0_avalon_slave_address),             //                          Timer_64Bit_0_avalon_slave.address
		.Timer_64Bit_0_avalon_slave_write                          (mm_interconnect_0_timer_64bit_0_avalon_slave_write),               //                                                    .write
		.Timer_64Bit_0_avalon_slave_read                           (mm_interconnect_0_timer_64bit_0_avalon_slave_read),                //                                                    .read
		.Timer_64Bit_0_avalon_slave_readdata                       (mm_interconnect_0_timer_64bit_0_avalon_slave_readdata),            //                                                    .readdata
		.Timer_64Bit_0_avalon_slave_writedata                      (mm_interconnect_0_timer_64bit_0_avalon_slave_writedata),           //                                                    .writedata
		.usb_gpx_s1_address                                        (mm_interconnect_0_usb_gpx_s1_address),                             //                                          usb_gpx_s1.address
		.usb_gpx_s1_readdata                                       (mm_interconnect_0_usb_gpx_s1_readdata),                            //                                                    .readdata
		.usb_irq_s1_address                                        (mm_interconnect_0_usb_irq_s1_address),                             //                                          usb_irq_s1.address
		.usb_irq_s1_readdata                                       (mm_interconnect_0_usb_irq_s1_readdata),                            //                                                    .readdata
		.usb_rst_s1_address                                        (mm_interconnect_0_usb_rst_s1_address),                             //                                          usb_rst_s1.address
		.usb_rst_s1_write                                          (mm_interconnect_0_usb_rst_s1_write),                               //                                                    .write
		.usb_rst_s1_readdata                                       (mm_interconnect_0_usb_rst_s1_readdata),                            //                                                    .readdata
		.usb_rst_s1_writedata                                      (mm_interconnect_0_usb_rst_s1_writedata),                           //                                                    .writedata
		.usb_rst_s1_chipselect                                     (mm_interconnect_0_usb_rst_s1_chipselect),                          //                                                    .chipselect
		.vga_display_0_avalon_slave_address                        (mm_interconnect_0_vga_display_0_avalon_slave_address),             //                          vga_display_0_avalon_slave.address
		.vga_display_0_avalon_slave_write                          (mm_interconnect_0_vga_display_0_avalon_slave_write),               //                                                    .write
		.vga_display_0_avalon_slave_read                           (mm_interconnect_0_vga_display_0_avalon_slave_read),                //                                                    .read
		.vga_display_0_avalon_slave_readdata                       (mm_interconnect_0_vga_display_0_avalon_slave_readdata),            //                                                    .readdata
		.vga_display_0_avalon_slave_writedata                      (mm_interconnect_0_vga_display_0_avalon_slave_writedata)            //                                                    .writedata
	);

	soc_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (pll_c0_clk),                             //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_c2_clk),                         //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
