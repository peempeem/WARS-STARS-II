	component soc is
		port (
			clk_clk             : in    std_logic                     := 'X';             -- clk
			reset_reset_n       : in    std_logic                     := 'X';             -- reset_n
			sdram_clk_clk       : out   std_logic;                                        -- clk
			sdram_wire_addr     : out   std_logic_vector(12 downto 0);                    -- addr
			sdram_wire_ba       : out   std_logic_vector(1 downto 0);                     -- ba
			sdram_wire_cas_n    : out   std_logic;                                        -- cas_n
			sdram_wire_cke      : out   std_logic;                                        -- cke
			sdram_wire_cs_n     : out   std_logic;                                        -- cs_n
			sdram_wire_dq       : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
			sdram_wire_dqm      : out   std_logic_vector(1 downto 0);                     -- dqm
			sdram_wire_ras_n    : out   std_logic;                                        -- ras_n
			sdram_wire_we_n     : out   std_logic;                                        -- we_n
			spi0_MISO           : in    std_logic                     := 'X';             -- MISO
			spi0_MOSI           : out   std_logic;                                        -- MOSI
			spi0_SCLK           : out   std_logic;                                        -- SCLK
			spi0_SS_n           : out   std_logic;                                        -- SS_n
			usb_gpx_export      : in    std_logic                     := 'X';             -- export
			usb_irq_export      : in    std_logic                     := 'X';             -- export
			usb_rst_export      : out   std_logic;                                        -- export
			vga_port_blue       : out   std_logic_vector(3 downto 0);                     -- blue
			vga_port_green      : out   std_logic_vector(3 downto 0);                     -- green
			vga_port_hs         : out   std_logic;                                        -- hs
			vga_port_red        : out   std_logic_vector(3 downto 0);                     -- red
			vga_port_vs         : out   std_logic;                                        -- vs
			i2c_conduit_data_in : in    std_logic                     := 'X';             -- conduit_data_in
			i2c_conduit_clk_in  : in    std_logic                     := 'X';             -- conduit_clk_in
			i2c_conduit_data_oe : out   std_logic;                                        -- conduit_data_oe
			i2c_conduit_clk_oe  : out   std_logic                                         -- conduit_clk_oe
		);
	end component soc;

	u0 : component soc
		port map (
			clk_clk             => CONNECTED_TO_clk_clk,             --        clk.clk
			reset_reset_n       => CONNECTED_TO_reset_reset_n,       --      reset.reset_n
			sdram_clk_clk       => CONNECTED_TO_sdram_clk_clk,       --  sdram_clk.clk
			sdram_wire_addr     => CONNECTED_TO_sdram_wire_addr,     -- sdram_wire.addr
			sdram_wire_ba       => CONNECTED_TO_sdram_wire_ba,       --           .ba
			sdram_wire_cas_n    => CONNECTED_TO_sdram_wire_cas_n,    --           .cas_n
			sdram_wire_cke      => CONNECTED_TO_sdram_wire_cke,      --           .cke
			sdram_wire_cs_n     => CONNECTED_TO_sdram_wire_cs_n,     --           .cs_n
			sdram_wire_dq       => CONNECTED_TO_sdram_wire_dq,       --           .dq
			sdram_wire_dqm      => CONNECTED_TO_sdram_wire_dqm,      --           .dqm
			sdram_wire_ras_n    => CONNECTED_TO_sdram_wire_ras_n,    --           .ras_n
			sdram_wire_we_n     => CONNECTED_TO_sdram_wire_we_n,     --           .we_n
			spi0_MISO           => CONNECTED_TO_spi0_MISO,           --       spi0.MISO
			spi0_MOSI           => CONNECTED_TO_spi0_MOSI,           --           .MOSI
			spi0_SCLK           => CONNECTED_TO_spi0_SCLK,           --           .SCLK
			spi0_SS_n           => CONNECTED_TO_spi0_SS_n,           --           .SS_n
			usb_gpx_export      => CONNECTED_TO_usb_gpx_export,      --    usb_gpx.export
			usb_irq_export      => CONNECTED_TO_usb_irq_export,      --    usb_irq.export
			usb_rst_export      => CONNECTED_TO_usb_rst_export,      --    usb_rst.export
			vga_port_blue       => CONNECTED_TO_vga_port_blue,       --   vga_port.blue
			vga_port_green      => CONNECTED_TO_vga_port_green,      --           .green
			vga_port_hs         => CONNECTED_TO_vga_port_hs,         --           .hs
			vga_port_red        => CONNECTED_TO_vga_port_red,        --           .red
			vga_port_vs         => CONNECTED_TO_vga_port_vs,         --           .vs
			i2c_conduit_data_in => CONNECTED_TO_i2c_conduit_data_in, --        i2c.conduit_data_in
			i2c_conduit_clk_in  => CONNECTED_TO_i2c_conduit_clk_in,  --           .conduit_clk_in
			i2c_conduit_data_oe => CONNECTED_TO_i2c_conduit_data_oe, --           .conduit_data_oe
			i2c_conduit_clk_oe  => CONNECTED_TO_i2c_conduit_clk_oe   --           .conduit_clk_oe
		);

