/*
module i2s (
	input logic           clk,
                         reset
)

end module
/*
assign i2c_serial_ARDUINO_IO[15]_in = arduino_adc_ARDUINO_IO[15];
assign arduino_ado_ARDUINO_IO[15] = i2c_serial_ARDUINO_IO[15]_oe ? 1'b0 : 1 'bz;

assign i2c_serial_ARDUINO_IO[14]_in = arduino_adc_ARDUINO_IO[14];
assign arduino_adc_ARDUINO_IO[14] = i2c_serial_ARDUINO_IO[14]_oe ? 1'b0 : 1'bz;
*/